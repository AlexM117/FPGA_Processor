//Alex Marlow & Graham Boyer TCES 330

//hex decoder module
module HexaHex( Hex, C);


input [3:0] C;  //input for hex
output reg [0:6] Hex;  //output for all figure segments

always@( C) begin

//cases for output based on input C
 case(C)
     4'b0000 : Hex = 7'b0000001; //0
	  4'b0001 : Hex = 7'b1001111; //1
	  4'b0010 : Hex = 7'b0010010; //2
	  4'b0011 : Hex = 7'b0000110; //3
	  4'b0100 : Hex = 7'b1001100; //4
	  4'b0101 : Hex = 7'b0100100; //5
	  4'b0110 : Hex = 7'b0100000; //6
	  4'b0111 : Hex = 7'b0001111; //7
	  4'b1000 : Hex = 7'b0000000; //8
	  4'b1001 : Hex = 7'b0001100; //9
	  4'b1010 : Hex = 7'b0001000; //A
	  4'b1011 : Hex = 7'b1100000; //B
	  4'b1100 : Hex = 7'b0110001; //C
	  4'b1101 : Hex = 7'b1000010; //D
	  4'b1110 : Hex = 7'b0110000; //E
	  4'b1111 : Hex = 7'b0111000; //F
 endcase

end

endmodule 